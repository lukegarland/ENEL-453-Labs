library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


entity Lab5 is
port(
		clk 			: in 	std_logic;
		reset			: in 	std_logic;
		AM_FM_Select	: in 	std_logic;
		R2R_Output		: out 	std_logic_vector(4 downto 0);
);
end Lab5;


architecture Behaviour of Lab5 is 




begin



end Behaviour;


