library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity sine_LUT is 

Port (
		reset			: in std_logic;
		value_in 		: in std_logic_vector(15 downto 0);
		sine_value		: out std_logic_vector(5 downto 0)

);

end sine_LUT;

architecture Behaviour of sine_LUT is 


type waveform_LUT is array (0 to 65535) of integer;

constant SINE_array_5 : waveform_LUT := ((0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (16), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-16), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0)
);
constant Sine_array_6 : waveform_LUT :=( (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (32), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (31), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (30), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (29), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (28), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (27), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (26), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (25), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (24), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (23), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (22), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (21), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (20), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (19), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (18), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (17), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (16), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (15), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (14), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (13), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (12), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (11), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (10), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (9), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (8), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (7), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (6), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (5), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (4), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (3), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (2), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-32), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-31), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-30), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-29), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-28), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-27), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-26), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-25), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-24), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-23), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-22), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-21), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-20), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-19), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-18), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-17), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-16), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-15), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-14), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-13), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-12), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-11), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-10), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-9), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-8), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-7), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-6), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-5), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-4), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-3), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-2), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (-1), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0)
);

begin

	process(reset, value_in)
	begin

	if(reset = '1') then
		sine_value <= (others => '0');
	else
		sine_value		<= std_logic_vector(to_signed(SINE_array_6(to_integer(unsigned(value_in))),SINE_value'length));
	end if;
	
	end process;





end Behaviour;
