library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity wave_LUTs is 

Port (
		reset			: in std_logic;
		value_in 		: in std_logic_vector(8 downto 0);
		wave_select		: in std_logic_vector(1 downto 0);
		wave_value		: out std_logic_vector(8 downto 0)

);

end wave_LUTs;


architecture Behaviour of wave_LUTs is 

component Mux4to1 is
	Generic ( busWidth : integer := 9); -- number to count       
	port(
	 selectLine : in std_logic_vector(1 downto 0);
	 input1 : in std_logic_vector(busWidth - 1 downto 0);
	 input2 : in std_logic_vector(busWidth - 1 downto 0);
	 input3 : in std_logic_vector(busWidth - 1 downto 0);
	 input4 : in std_logic_vector(busWidth - 1 downto 0);
	 muxOutput : out std_logic_vector(busWidth - 1 downto 0)
	 );
end component;


type waveform_LUT is array (0 to 511) of integer;

constant SQUARE_LUT : waveform_LUT := (
(0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (0), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1), (1)
);
constant SAWTOOTH_LUT : waveform_LUT := (
(0), (1), (2), (3), (4), (5), (6), (7), (8), (9), (10), (11), (12), (13), (14), (15), (16), (17), (18), (19), (20), (21), (22), (23), (24), (25), (26), (27), (28), (29), (30), (31), (32), (33), (34), (35), (36), (37), (38), (39), (40), (41), (42), (43), (44), (45), (46), (47), (48), (49), (50), (51), (52), (53), (54), (55), (56), (57), (58), (59), (60), (61), (62), (63), (64), (65), (66), (67), (68), (69), (70), (71), (72), (73), (74), (75), (76), (77), (78), (79), (80), (81), (82), (83), (84), (85), (86), (87), (88), (89), (90), (91), (92), (93), (94), (95), (96), (97), (98), (99), (100), (101), (102), (103), (104), (105), (106), (107), (108), (109), (110), (111), (112), (113), (114), (115), (116), (117), (118), (119), (120), (121), (122), (123), (124), (125), (126), (127), (128), (129), (130), (131), (132), (133), (134), (135), (136), (137), (138), (139), (140), (141), (142), (143), (144), (145), (146), (147), (148), (149), (150), (151), (152), (153), (154), (155), (156), (157), (158), (159), (160), (161), (162), (163), (164), (165), (166), (167), (168), (169), (170), (171), (172), (173), (174), (175), (176), (177), (178), (179), (180), (181), (182), (183), (184), (185), (186), (187), (188), (189), (190), (191), (192), (193), (194), (195), (196), (197), (198), (199), (200), (201), (202), (203), (204), (205), (206), (207), (208), (209), (210), (211), (212), (213), (214), (215), (216), (217), (218), (219), (220), (221), (222), (223), (224), (225), (226), (227), (228), (229), (230), (231), (232), (233), (234), (235), (236), (237), (238), (239), (240), (241), (242), (243), (244), (245), (246), (247), (248), (249), (250), (251), (252), (253), (254), (255), (256), (257), (258), (259), (260), (261), (262), (263), (264), (265), (266), (267), (268), (269), (270), (271), (272), (273), (274), (275), (276), (277), (278), (279), (280), (281), (282), (283), (284), (285), (286), (287), (288), (289), (290), (291), (292), (293), (294), (295), (296), (297), (298), (299), (300), (301), (302), (303), (304), (305), (306), (307), (308), (309), (310), (311), (312), (313), (314), (315), (316), (317), (318), (319), (320), (321), (322), (323), (324), (325), (326), (327), (328), (329), (330), (331), (332), (333), (334), (335), (336), (337), (338), (339), (340), (341), (342), (343), (344), (345), (346), (347), (348), (349), (350), (351), (352), (353), (354), (355), (356), (357), (358), (359), (360), (361), (362), (363), (364), (365), (366), (367), (368), (369), (370), (371), (372), (373), (374), (375), (376), (377), (378), (379), (380), (381), (382), (383), (384), (385), (386), (387), (388), (389), (390), (391), (392), (393), (394), (395), (396), (397), (398), (399), (400), (401), (402), (403), (404), (405), (406), (407), (408), (409), (410), (411), (412), (413), (414), (415), (416), (417), (418), (419), (420), (421), (422), (423), (424), (425), (426), (427), (428), (429), (430), (431), (432), (433), (434), (435), (436), (437), (438), (439), (440), (441), (442), (443), (444), (445), (446), (447), (448), (449), (450), (451), (452), (453), (454), (455), (456), (457), (458), (459), (460), (461), (462), (463), (464), (465), (466), (467), (468), (469), (470), (471), (472), (473), (474), (475), (476), (477), (478), (479), (480), (481), (482), (483), (484), (485), (486), (487), (488), (489), (490), (491), (492), (493), (494), (495), (496), (497), (498), (499), (500), (501), (502), (503), (504), (505), (506), (507), (508), (509), (510), (511)
);

constant TRIANGLE_LUT : waveform_LUT := (
(0), (2), (4), (6), (8), (10), (12), (14), (16), (18), (20), (22), (24), (26), (28), (30), (32), (34), (36), (38), (40), (42), (44), (46), (48), (50), (52), (54), (56), (58), (60), (62), (64), (66), (68), (70), (72), (74), (76), (78), (80), (82), (84), (86), (88), (90), (92), (94), (96), (98), (100), (102), (104), (106), (108), (110), (112), (114), (116), (118), (120), (122), (124), (126), (128), (130), (132), (134), (136), (138), (140), (142), (144), (146), (148), (150), (152), (154), (156), (158), (160), (162), (164), (166), (168), (170), (172), (174), (176), (178), (180), (182), (184), (186), (188), (190), (192), (194), (196), (198), (200), (202), (204), (206), (208), (210), (212), (214), (216), (218), (220), (222), (224), (226), (228), (230), (232), (234), (236), (238), (240), (242), (244), (246), (248), (250), (252), (254), (256), (258), (260), (262), (264), (266), (268), (270), (272), (274), (276), (278), (280), (282), (284), (286), (288), (290), (292), (294), (296), (298), (300), (302), (304), (306), (308), (310), (312), (314), (316), (318), (320), (322), (324), (326), (328), (330), (332), (334), (336), (338), (340), (342), (344), (346), (348), (350), (352), (354), (356), (358), (360), (362), (364), (366), (368), (370), (372), (374), (376), (378), (380), (382), (384), (386), (388), (390), (392), (394), (396), (398), (400), (402), (404), (406), (408), (410), (412), (414), (416), (418), (420), (422), (424), (426), (428), (430), (432), (434), (436), (438), (440), (442), (444), (446), (448), (450), (452), (454), (456), (458), (460), (462), (464), (466), (468), (470), (472), (474), (476), (478), (480), (482), (484), (486), (488), (490), (492), (494), (496), (498), (500), (502), (504), (506), (508), (510), (510), (508), (506), (504), (502), (500), (498), (496), (494), (492), (490), (488), (486), (484), (482), (480), (478), (476), (474), (472), (470), (468), (466), (464), (462), (460), (458), (456), (454), (452), (450), (448), (446), (444), (442), (440), (438), (436), (434), (432), (430), (428), (426), (424), (422), (420), (418), (416), (414), (412), (410), (408), (406), (404), (402), (400), (398), (396), (394), (392), (390), (388), (386), (384), (382), (380), (378), (376), (374), (372), (370), (368), (366), (364), (362), (360), (358), (356), (354), (352), (350), (348), (346), (344), (342), (340), (338), (336), (334), (332), (330), (328), (326), (324), (322), (320), (318), (316), (314), (312), (310), (308), (306), (304), (302), (300), (298), (296), (294), (292), (290), (288), (286), (284), (282), (280), (278), (276), (274), (272), (270), (268), (266), (264), (262), (260), (258), (256), (254), (252), (250), (248), (246), (244), (242), (240), (238), (236), (234), (232), (230), (228), (226), (224), (222), (220), (218), (216), (214), (212), (210), (208), (206), (204), (202), (200), (198), (196), (194), (192), (190), (188), (186), (184), (182), (180), (178), (176), (174), (172), (170), (168), (166), (164), (162), (160), (158), (156), (154), (152), (150), (148), (146), (144), (142), (140), (138), (136), (134), (132), (130), (128), (126), (124), (122), (120), (118), (116), (114), (112), (110), (108), (106), (104), (102), (100), (98), (96), (94), (92), (90), (88), (86), (84), (82), (80), (78), (76), (74), (72), (70), (68), (66), (64), (62), (60), (58), (56), (54), (52), (50), (48), (46), (44), (42), (40), (38), (36), (34), (32), (30), (28), (26), (24), (22), (20), (18), (16), (14), (12), (10), (8), (6), (4), (2), (0)
);

constant SINE_LUT : waveform_LUT := (
(256), (259), (262), (265), (268), (271), (274), (277), (280), (284), (287), (290), (293), (296), (299), (302), (305), (308), (311), (314), (317), (320), (324), (327), (330), (333), (335), (338), (341), (344), (347), (350), (353), (356), (359), (362), (365), (367), (370), (373), (376), (378), (381), (384), (387), (389), (392), (395), (397), (400), (402), (405), (407), (410), (412), (415), (417), (420), (422), (424), (427), (429), (431), (434), (436), (438), (440), (442), (444), (447), (449), (451), (453), (455), (457), (458), (460), (462), (464), (466), (468), (469), (471), (473), (474), (476), (477), (479), (480), (482), (483), (485), (486), (487), (489), (490), (491), (492), (493), (495), (496), (497), (498), (499), (500), (500), (501), (502), (503), (504), (504), (505), (506), (506), (507), (507), (508), (508), (509), (509), (509), (510), (510), (510), (510), (510), (510), (510), (511), (510), (510), (510), (510), (510), (510), (510), (509), (509), (509), (508), (508), (507), (507), (506), (506), (505), (504), (504), (503), (502), (501), (500), (500), (499), (498), (497), (496), (495), (493), (492), (491), (490), (489), (487), (486), (485), (483), (482), (480), (479), (477), (476), (474), (473), (471), (469), (468), (466), (464), (462), (460), (458), (457), (455), (453), (451), (449), (447), (444), (442), (440), (438), (436), (434), (431), (429), (427), (424), (422), (420), (417), (415), (412), (410), (407), (405), (402), (400), (397), (395), (392), (389), (387), (384), (381), (378), (376), (373), (370), (367), (365), (362), (359), (356), (353), (350), (347), (344), (341), (338), (335), (333), (330), (327), (324), (320), (317), (314), (311), (308), (305), (302), (299), (296), (293), (290), (287), (284), (280), (277), (274), (271), (268), (265), (262), (259), (256), (253), (250), (247), (244), (241), (238), (235), (232), (228), (225), (222), (219), (216), (213), (210), (207), (204), (201), (198), (195), (192), (188), (185), (182), (179), (177), (174), (171), (168), (165), (162), (159), (156), (153), (150), (147), (145), (142), (139), (136), (134), (131), (128), (125), (123), (120), (117), (115), (112), (110), (107), (105), (102), (100), (97), (95), (92), (90), (88), (85), (83), (81), (78), (76), (74), (72), (70), (68), (65), (63), (61), (59), (57), (55), (54), (52), (50), (48), (46), (44), (43), (41), (39), (38), (36), (35), (33), (32), (30), (29), (27), (26), (25), (23), (22), (21), (20), (19), (17), (16), (15), (14), (13), (12), (12), (11), (10), (9), (8), (8), (7), (6), (6), (5), (5), (4), (4), (3), (3), (3), (2), (2), (2), (2), (2), (2), (2), (1), (2), (2), (2), (2), (2), (2), (2), (3), (3), (3), (4), (4), (5), (5), (6), (6), (7), (8), (8), (9), (10), (11), (12), (12), (13), (14), (15), (16), (17), (19), (20), (21), (22), (23), (25), (26), (27), (29), (30), (32), (33), (35), (36), (38), (39), (41), (43), (44), (46), (48), (50), (52), (54), (55), (57), (59), (61), (63), (65), (68), (70), (72), (74), (76), (78), (81), (83), (85), (88), (90), (92), (95), (97), (100), (102), (105), (107), (110), (112), (115), (117), (120), (123), (125), (128), (131), (134), (136), (139), (142), (145), (147), (150), (153), (156), (159), (162), (165), (168), (171), (174), (177), (179), (182), (185), (188), (192), (195), (198), (201), (204), (207), (210), (213), (216), (219), (222), (225), (228), (232), (235), (238), (241), (244), (247), (250), (253)
);

signal SQUARE_value: std_logic_vector(8 downto 0);
signal SAWTOOTH_value:  std_logic_vector(8 downto 0);
signal TRIANGLE_value:  std_logic_vector(8 downto 0);
signal SINE_value:  std_logic_vector(8 downto 0);
signal wave_value_from_mux:  std_logic_vector(8 downto 0);




begin

	process(reset, value_in, wave_select)
	begin

	if(reset = '1') then
		wave_value <= (others => '0');
	else
		wave_value 		<= wave_value_from_mux;
	end if;
	
	end process;
	
	
		SQUARE_value 	<= std_logic_vector(to_unsigned(SQUARE_LUT(to_integer(unsigned(value_in))),SQUARE_value'length));
		SAWTOOTH_value 	<= std_logic_vector(to_unsigned(SAWTOOTH_LUT(to_integer(unsigned(value_in))),SAWTOOTH_value'length));
		TRIANGLE_value 	<= std_logic_vector(to_unsigned(TRIANGLE_LUT(to_integer(unsigned(value_in))),TRIANGLE_value'length));
		SINE_value		<= std_logic_vector(to_unsigned(SINE_LUT(to_integer(unsigned(value_in))),SINE_value'length));
	Select_wave_ins: Mux4to1
					generic map (busWidth => 9)
					port map(
						selectLine	=> wave_select,
						input1 		=> SQUARE_value,
						input2		=> SAWTOOTH_value,
						input3		=> TRIANGLE_value,
						input4		=> SINE_value,
						muxOutput	=> wave_value_from_mux
					);



end Behaviour;
